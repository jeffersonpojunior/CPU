module control_unit(); // Mini CPU