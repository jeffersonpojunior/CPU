module memory();