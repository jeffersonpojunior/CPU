module alu(); // Arithmetic logic unit